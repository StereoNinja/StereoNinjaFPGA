module Ram_Controller(input write_read_n,clk,reset,input[7:0] red)
		
		
end module;